`timescale 1ns/1ps

module permitation_xor import ascon_pack::*;
   (
    input logic 	clock_i,
    input logic 	resetb_i,
    input logic 	select_i,
    input 		type_state permutation_i,
    input logic [3:0] 	roundp_i,
    input logic [63:0] 	data_xor_up_i,
    input logic [255:0] data_xor_down_i,
    input logic 	ena_xor_up_i,
    input logic 	ena_xor_down_i,
    input logic 	ena_reg_i,
    output 		type_state permutation_o,
    output type_state  xor_up_o
    );

   //selection de l'entree par un multiplexeur
   type_state state_mux;
   assign state_mux = (select_i) ? permutation_i : permutation_o;

   //xor up et nultiplexeur pour selectionner l'entree
   type_state state_pc;
   assign state_pc[0] = (ena_xor_up_i==1'b1) ? state_mux[0]^data_xor_up_i : state_mux[0];
   assign state_pc[1] = state_mux[1];
   assign state_pc[2] = state_mux[2];
   assign state_pc[3] = state_mux[3];
   assign state_pc[4] = state_mux[4];

  
   type_state state_ps;
   //permutation constante
   permitation_constante pc(
			    .constante_add_i(state_pc),
			    .round_i(roundp_i),
			    .constante_add_o(state_ps)
			    );

   type_state state_pl;
   //permutation de substitution
   permitation_substitution ps(
			       .substitution_i(state_ps),
			       .substitution_o(state_pl)
			       );
   type_state state_p;
   //permutation de diffusion lineaire
   permitation_diffusion pl(
			    .diffusion_i(state_pl),
			    .diffusion_o(state_p)
			    );

   //xor down et multiplexeur pour choisir la sortie
    type_state state_mux_p;
   assign state_mux_p[0] = state_p[0];
   assign state_mux_p[1] = (ena_xor_down_i==1'b1) ? state_p[1]^data_xor_down_i[255:192] : state_p[1];
   assign state_mux_p[2] = (ena_xor_down_i==1'b1) ? state_p[2]^data_xor_down_i[191:128] : state_p[2];
   assign state_mux_p[3] = (ena_xor_down_i==1'b1) ? state_p[3]^data_xor_down_i[127:64] : state_p[3];
   assign state_mux_p[4] = (ena_xor_down_i==1'b1) ? state_p[4]^data_xor_down_i[63:0] : state_p[4];

   //registre de memorisation
   always @ (posedge clock_i, negedge resetb_i) begin
      if(resetb_i == 1'b0) begin
	 permutation_o <= {64'h0,64'h0,64'h0,64'h0,64'h0};
      end
      else begin
	 if(ena_reg_i==1'b1)begin 
            permutation_o <= state_mux_p;
	 end
      end
   end

   assign xor_up_o = state_pc;
endmodule : permitation_xor
